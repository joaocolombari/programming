--
--

package riscv_pkg is


end package;


package body riscv_pkg is


end package body;